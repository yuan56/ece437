mg252@cparch06.ecn.purdue.edu.17839:1422840629