mg252@cparch03.ecn.purdue.edu.9362:1422840637